

module data_maker(
    output wire [31:0] data1,
    output wire [31:0] data2,
    output wire [31:0] data3,
    output wire [31:0] data4
    );

assign data1 = 32'd520;
assign data2 = 32'd778;
assign data3 = 32'd2022;
assign data4 = 32'd1234;
    
endmodule
